import lc3b_types::*;

module fetch_logic
(
    input lc3b_mem_wmask in,
	 output lc3b_mux_sel out
);

always_comb
begin

end

endmodule : fetch_logic
