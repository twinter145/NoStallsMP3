import lc3b_types::*;

module datapath
(
	/* inputs */
	input clk,
	
	/* outputs */
);
//internal signals


//fetch


//decode


//execute


//memory


//write back


endmodule : datapath
